library verilog;
use verilog.vl_types.all;
entity operator_adapter_vlg_vec_tst is
end operator_adapter_vlg_vec_tst;
