library verilog;
use verilog.vl_types.all;
entity arithmetic_vlg_vec_tst is
end arithmetic_vlg_vec_tst;
