library verilog;
use verilog.vl_types.all;
entity divider_vlg_vec_tst is
end divider_vlg_vec_tst;
