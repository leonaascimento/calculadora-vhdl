library verilog;
use verilog.vl_types.all;
entity subtractor_vlg_vec_tst is
end subtractor_vlg_vec_tst;
