library verilog;
use verilog.vl_types.all;
entity pwm_controller_vlg_vec_tst is
end pwm_controller_vlg_vec_tst;
