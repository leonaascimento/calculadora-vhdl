library verilog;
use verilog.vl_types.all;
entity pwm_module_vlg_vec_tst is
end pwm_module_vlg_vec_tst;
